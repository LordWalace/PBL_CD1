//module matriz(Alto, Medio, Baixo, D1, D2, D3, A7, B7, C7, D7, E7, F7, G7);
	
//	input Alto, Medio, Baixo;
//	output 

//endmodule 